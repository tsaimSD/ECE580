module no_branch_predictor;
  // This is a placeholder module to avoid elaboration errors.
  // It contains no logic because we assume NO branch prediction in this model.
endmodule